
-- synthesis translate_on
architecture rtl of fifo is

-- synopsis something
  alias designator is name;

-- Random comment
  alias designator is name;

-- altera something
  alias designator is name;

-- xilinx something

begin
-- RTL_SYNTHESIS ON
end architecture rtl;
-- synthesis translate_off
